module helloV;
    initial
    begin
        $display("Learning something new today");
        $display("Yes, Hello World HDL");
    end
endmodule
